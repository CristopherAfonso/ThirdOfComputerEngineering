library verilog;
use verilog.vl_types.all;
entity pr1_cpu_extendida is
end pr1_cpu_extendida;
